module v2

#pkgconfig gio-2.0
#flag -Wno-deprecated-declarations
